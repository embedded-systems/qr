#include "connection_builder.vh"

#bigfunc ADD_1TO1_INPUT_DEVICE(NAME, INDEX, INT_INDX, WIDTH, PINS)
	REGISTER_INPUT_PIN(NAME, WIDTH, PINS)
	CREATE_MUX_ENTRY(INDEX, NAME, WIDTH, NAME, '1')
	CREATE_INTERRUPT_ON_CHANGE(INT_INDX, NAME, WIDTH)
#endbigfunc

#bigfunc ADD_1TO1_OUTPUT_DEVICE(NAME, INDEX, WIDTH, PINS)
	REGISTER_OUTPUT_PIN(NAME, WIDTH, PINS)
	CREATE_REGISTER(INDEX, NAME_reg, WIDTH, NAME)
	#ifdef __IN_VHDL 
		NAME <= NAME_reg;
	#endif 
#endbigfunc

