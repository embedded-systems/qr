-------------------------------------------------------------------------------
-- Filename:             sram-32.vhd
-- Entity:               sram32
-- Architectures:        behaviour
-- Author:               Sijmen Woutersen
-- Last Modified:        2007/01/06
-- Version:              1.0
-- Description:          Memory controller for the X32 on the spartan 3 starter
--                       board. The memory controller transforms X32 memory
--                       operations into operations supported by the memory 
--                       chips of the board. A decoder is used to decode the
--                       unaligned data into aligned data (and visa versa), as
--                       the memory chips require data to be aligned, while the
--                       X32 reads from/writes to unlaligned addresses
--
-- 	Copyright (c) 2005-2007, Software Technology Department, TU Delft
--	All rights reserved.
--
-- 	This program is free software; you can redistribute it and/or
--	modify it under the terms of the GNU General Public License
--	as published by the Free Software Foundation; either version 2
--	of the License, or (at your option) any later version.
--	
--	This program is distributed in the hope that it will be useful,
-- 	but WITHOUT ANY WARRANTY; without even the implied warranty of
--	MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--	GNU General Public License for more details.
--	
--	You should have received a copy of the GNU General Public License
--	along with this program; if not, write to the Free Software
-- 	Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA  
--  02111-1307, USA.
--	
--  See the GNU General Public License here:
--
--  http://www.gnu.org/copyleft/gpl.html#SEC1
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.types.all;

entity sram32 is
	port (
		-- system clock
		clk							: in    std_logic;
		-- system reset
		reset						: in    std_logic;
		
		-- memory address (unaligned)
		mem_address			: in    std_logic_vector(19 downto 0);
		-- data to memory
		mem_data_in			: in    std_logic_vector(31 downto 0);
		-- data from memory
		mem_data_out  	: out   std_logic_vector(31 downto 0);
		-- size of data (see types.vhd)
		mem_data_size		: in    std_logic_vector(2 downto 0);
		-- data signedness (1=signed, 0=unsigned)
		mem_data_signed	: in    std_logic;
		-- start read operation (high = start read)
		mem_read				: in    std_logic;
		-- start write operation (high = start write)
		mem_write				: in    std_logic;
		-- pulses high when the operation finishes
		mem_ready				: out   std_logic;

		-- sram address (32-bit aligned, both chips)
		sram_address		: out   std_logic_vector(17 downto 0);
		-- chip enable (chip 1)
		sram_ce1				: out   std_logic;
		-- upper byte enable (chip 1)
		sram_ub1				: out   std_logic;
		-- lower byte enable (chip 1)
		sram_lb1				: out   std_logic;
		-- memory data (chip 1)
		sram_data1			: inout std_logic_vector(15 downto 0);
		-- chip enable (chip 2)
		sram_ce2				: out   std_logic;
		-- upper byte enable (chip 2)
		sram_ub2				: out   std_logic;
		-- lower byte enable (chip 2)
		sram_lb2				: out   std_logic;
		-- memory data (chip 2)
		sram_data2			: inout std_logic_vector(15 downto 0);
		-- output enable (both chips)
		sram_oe					: out   std_logic;
		-- write enable (both chips)
		sram_we					: out   std_logic;

		-- overflow, as generated by the decoder
		overflow				: out	std_logic
	);
	
end entity;

architecture behaviour of sram32 is
	-- fsm states
	type STATE_TYPE is (RESET_STATE, IDLE, READ_WORD1B, 
		READ_WORD2A, READ_WORD2B, WRITE_WORD1, WRITE_WORD2, 
		ALIGN_OUTPUT_DATA, ALIGN_INPUT_DATA);
	signal state_i, state_o : STATE_TYPE;
	
	-- lower & upper aligned memory addresses:
	--  when address = 0x03, then mem_address1 = 0x00 and
	--  mem_address2 = 0x01, as when reading 32-bit, data
	--  from both addresses is required
	signal mem_address1 : std_logic_vector(17 downto 0);
	signal mem_address2 : std_logic_vector(17 downto 0);

	-- data signals
	signal mem_data_in1, mem_data_out1_i, mem_data_out2_i, 
		mem_data_out1_o, mem_data_out2_o : std_logic_vector(31 downto 0);
	signal mem_data_in2 : std_logic_vector(31 downto 8);
	
	-- byte enable signals
	signal bytes_enable1_i, bytes_enable2_i, bytes_enable1_o, bytes_enable2_o, 
		bytes_enable : std_logic_vector(3 downto 0);

	-- memory decoder (see mem_decoder.vhd)
	component mem_decoder is
		port (
			address_offset 	: in  std_logic_vector(1 downto 0);
			mem_data_size		: in  std_logic_vector(2 downto 0);
			mem_data_signed	: in  std_logic;
			
			mem_data_in1		: in  std_logic_vector(31 downto 0);
			mem_data_in2		: in  std_logic_vector(31 downto 8);
			proc_data_in		: out std_logic_vector(31 downto 0);
			
			proc_data_out		: in  std_logic_vector(31 downto 0);
			mem_data_out1		: out std_logic_vector(31 downto 0);
			mem_data_out2		: out std_logic_vector(31 downto 0);
			
			bytes_enable1		: out std_logic_vector(3 downto 0);
			bytes_enable2		: out std_logic_vector(3 downto 0);

			overflow		: out std_logic
		);
	end component;
	
	-- register store sginals
	signal store1, store2, store_addr, store_outputs : std_logic;

	signal mem_address_offset : std_logic_vector(1 downto 0);
	signal sig_overflow : std_logic;
begin
	-- overflow only on write
	overflow <= sig_overflow and mem_write;

	-- memory decoder
	dec: mem_decoder port map(mem_address_offset, mem_data_size, mem_data_signed,
		mem_data_in1, mem_data_in2, mem_data_out, mem_data_in, 
		mem_data_out1_i, mem_data_out2_i, bytes_enable1_i, bytes_enable2_i,
		sig_overflow);

	-- always enable both chips
	sram_ce1 <= '0';
	sram_ce2 <= '0';

	-- byte enable signals
	sram_ub1 <= bytes_enable(3);
	sram_lb1 <= bytes_enable(2);
	sram_ub2 <= bytes_enable(1);
	sram_lb2 <= bytes_enable(0);

	process(state_o, mem_read, mem_write, bytes_enable1_o, bytes_enable2_o, 
		mem_data_out1_o, mem_data_out2_o, mem_address1, mem_address2,
		bytes_enable2_i, mem_address) begin
		
		case state_o is
			when RESET_STATE =>
				-- reset/startup stage
				mem_ready <= '0';

				sram_data1 <= (others => '-');
				sram_data2 <= (others => '-');
				bytes_enable <= (others => '-');
				sram_address <= (others => '-');
				
				sram_we <= '1';
				sram_oe <= '1';
				
				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

				state_i <= IDLE;
			when IDLE =>
				-- idle, wait for read/write operations
				mem_ready <= '0';

				sram_data1 <= (others => '-');
				sram_data2 <= (others => '-');
				-- already enable all bytes, and read from the lower address,
				-- such that the first word is read immediatly when reading data
				bytes_enable <= "0000";
				sram_address <= mem_address(19 downto 2);

				-- output enable, but not write enable
				sram_we <= '1';
				sram_oe <= '0';

				-- store only the address+1, so that the high address is
				-- already available in the next state
				store1 <= '0';
				store2 <= '0';
				store_addr <= '1';
				store_outputs <= '0';
				
				if (mem_read = '1') then
					-- continue reading
					state_i <= READ_WORD1B;
				elsif (mem_write = '1') then
					-- TODO: can the compute outputs state be included in the idle state?
					state_i <= ALIGN_OUTPUT_DATA;
				else
					state_i <= IDLE;
				end if;
			-- THIS STATE IS NOW (MAY 11 2006) INCLUDED IN THE IDLE STATE
			--when READ_WORD1A =>
			--	mem_ready <= '0';

			--	sram_data1 <= (others => 'Z');
			--	sram_data2 <= (others => 'Z');
			--	bytes_enable <= "0000";
			--	sram_address <= mem_address1;

			--	sram_we <= '1';
			--	sram_oe <= '0';

			--	store1 <= '0';
			--	store2 <= '0';
			--	store_addr <= '0';
			--	store_outputs <= '0';

			--	state_i <= READ_WORD1B;
			when READ_WORD1B =>
				-- save word 1 from memory
				mem_ready <= '0';

				sram_data1 <= (others => 'Z');
				sram_data2 <= (others => 'Z');
				bytes_enable <= "0000";
				sram_address <= mem_address1;

				sram_we <= '1';
				sram_oe <= '0';

				store1 <= '1';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

				-- if only 1 word needs to be read, continue to alignment
				if (bytes_enable2_i = "1111") then
					state_i <= ALIGN_INPUT_DATA;
				else
					state_i <= READ_WORD2A;
				end if;
			when READ_WORD2A =>
				-- update memory signals to read word 2
				mem_ready <= '0';

				sram_data1 <= (others => 'Z');
				sram_data2 <= (others => 'Z');
				bytes_enable <= "0000";
				sram_address <= mem_address2;

				sram_we <= '1';
				sram_oe <= '0';

				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

				state_i <= READ_WORD2B;
			when READ_WORD2B =>
				-- save word 2
				mem_ready <= '0';

				sram_data1 <= (others => 'Z');
				sram_data2 <= (others => 'Z');
				bytes_enable <= "0000";
				sram_address <= mem_address2;

				sram_we <= '1';
				sram_oe <= '0';

				store1 <= '0';
				store2 <= '1';
				store_addr <= '0';
				store_outputs <= '0';

				state_i <= ALIGN_INPUT_DATA;
			when ALIGN_OUTPUT_DATA =>
				-- align the output data into two words
				mem_ready <= '0';

				sram_data1 <= (others => '-');
				sram_data2 <= (others => '-');
				bytes_enable <= (others => '-');
				sram_address <= (others => '-');
				
				sram_we <= '1';
				sram_oe <= '1';
				
				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '1';

				state_i <= WRITE_WORD1;
			when WRITE_WORD1 =>
				-- write word 1 
				--mem_ready <= '0';

				sram_data1 <= mem_data_out1_o(31 downto 16);
				sram_data2 <= mem_data_out1_o(15 downto 0);
				bytes_enable <= bytes_enable1_o;
				sram_address <= mem_address1;

				sram_we <= '0';
				sram_oe <= '1';

				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

				-- if only the lower word must be written, report ready
				if (bytes_enable2_i = "1111") then
					--state_i <= READY_STATE;
					state_i <= IDLE;
					mem_ready <= '1';
				else
					state_i <= WRITE_WORD2;
					mem_ready <= '0';
				end if;
			when WRITE_WORD2 =>
				-- write word 2
--				mem_ready <= '0';
				-- report ready
				mem_ready <= '1';

				sram_data1 <= mem_data_out2_o(31 downto 16);
				sram_data2 <= mem_data_out2_o(15 downto 0);
				bytes_enable <= bytes_enable2_o;
				sram_address <= mem_address2;

				sram_we <= '0';
				sram_oe <= '1';

				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

--				state_i <= READY_STATE;
				state_i <= IDLE;
--			when READY =>
			when ALIGN_INPUT_DATA =>
				-- align the 2 input words into a single word
				mem_ready <= '1';

				sram_we <= '1';
				sram_oe <= '1';

				sram_data1 <= (others => '-');
				sram_data2 <= (others => '-');
				bytes_enable <= (others => '-');
				sram_address <= (others => '-');

				store1 <= '0';
				store2 <= '0';
				store_addr <= '0';
				store_outputs <= '0';

				state_i <= IDLE;
		end case;
	end process;

	-- fsm register
	process(clk, reset, state_i) begin
		if (clk'event and clk = '1') then
			if (reset = '1') then
				state_o <= RESET_STATE;
			else
				state_o <= state_i;
			end if;
		end if;
	end process;

	-- (low) address register
	process(clk, reset, store_addr, mem_address) begin
		if (clk'event and clk = '1') then
			if (reset = '1') then
				mem_address1 <= (others => '0');
				mem_address_offset <= (others => '0');
			elsif (store_addr = '1') then
				mem_address1 <= mem_address(19 downto 2);
				mem_address_offset <= mem_address(1 downto 0);
			end if;
		end if;
	end process;	

	-- (high) address register
	process(clk, reset, mem_address1) begin
		if (clk'event and clk = '1') then
			if (reset = '1') then
				mem_address2 <= (others => '0');
			else
				mem_address2 <= mem_address1+1;
			end if;
		end if;
	end process;	

	-- low word register
	process(clk, reset, store1, mem_data_in1, sram_data1, sram_data2) begin
		if (clk'event and clk = '1') then
			if (reset = '1') then
				mem_data_in1 <= (others => '0');
			elsif (store1 = '1') then
				mem_data_in1(31 downto 16) <= sram_data1;
				mem_data_in1(15 downto 0) <= sram_data2;
			end if;
		end if;
	end process;	

	-- high word register
	process(clk, reset, store2, mem_data_in2, sram_data1, sram_data2) begin
		if (clk'event and clk = '1') then
			if (reset = '1') then
				mem_data_in2 <= (others => '0');
			elsif (store2 = '1') then
				mem_data_in2(31 downto 16) <= sram_data1;
				mem_data_in2(15 downto 8) <= sram_data2(15 downto 8);
			end if;
		end if;
	end process;	

	-- decoded data register
	process(clk, reset, store_outputs, 
		mem_data_out1_i, mem_data_out2_i, bytes_enable1_i, bytes_enable2_i,
		mem_data_out1_o, mem_data_out2_o, bytes_enable1_o, bytes_enable2_o) begin
	
		if (clk'event and clk = '1') then
			if (reset = '1') then
				mem_data_out1_o <= (others => '0');
				mem_data_out2_o <= (others => '0');
				bytes_enable1_o <= (others => '0');
				bytes_enable2_o <= (others => '0');
			elsif (store_outputs = '1') then
				mem_data_out1_o <= mem_data_out1_i;
				mem_data_out2_o <= mem_data_out2_i;
				bytes_enable1_o <= bytes_enable1_i;
				bytes_enable2_o <= bytes_enable2_i;
			end if;
		end if;
	end process;	
	


end architecture;
